/**************************************************************************/
// Copyright (c) 2024, OASIS Lab
// MODULE: TETRIS
// FILE NAME: TETRIS_encrypted.v
// VERSRION: 1.0
// DATE: August 15, 2024
// AUTHOR: Yu-Hsuan Hsu, NYCU IEE
// DESCRIPTION: ICLAB2024FALL / LAB3 / TETRIS_demo
// MODIFICATION HISTORY:
// Date                 Description
// 
/**************************************************************************/
module TETRIS
`protected
gOF=^2&42fF#^Xgf:=-ZRBI933\4G2(,&])S+,F0.20[U)BQ)EH<,)+0HR@4XCZU
/H^Bf>3;+/0,>#0P+R=@B\[:B:9<[4NZ(bcdQ@098D<7f-H-5>bJ^cK#(a&==]cF
,Vf]5FJ3725AY[Q/g7-@VX[C(FFH:@=XbN(\V->R;8GFGQgQJAVHI]e<J\a7WJ>9
eQTXDE>OZNW-YgbZ_.O+AMBZ1U-S[T;?fG6HMGF__[.Hee?W67^Y29dPgLecI5+G
Ubf.dBB#e>8=/-P,;BB>9SEKc<>LDR@/+?[b00ZL,6F7G+U?.OK--b02495Ef9^=
9;ZJK,BHb\ZRVK,b;=^ZA-WgGF7XA)S@fQ+3&_2WI+]1>AfaSVC^D/BV?S6c5[2G
a^9BC5be#A>eB+<L0PW:Lf]#&OV6ebJE7O<+gWAD?5b#=3ZdUD9V3,AUKK[gW@JT
]aQXC7[8KO1P_AOL1^aD(VdKBc,Z.-FA:5X?<_X[7bbB.GGe;L?c><39XQABV4E/
bbU>9La.V=.=W&#Ta7UcVe>KUE<Q10=7X@,)5Z90838G0C8T#F,SHBX[Z#[#_O)2
@93,KU-;M)Df=&5[_AB5VV&b4MXUM]AI5d]dQ?9;H\Z,_3dZP>:H/:V\JGJ]Y8&;
E80:Y=OQJ,Z(bBUF9a1YdM2CfTB4BM/75JGI?\4:;,6.ce2J.A64P+d79@XO8(UT
fS@]dC\C;4c/4O2RcY>8O=cL,O]NPN\,K@^D8<HV]T=8P/Dg?Y9e,(FG4P7]L>N7
PIX#QNU?F)&FOOE[3@AE@^R6H3M,S4ff^f2>@gcC^I?8[Pe&?@aOBR9)M7YfEAO:
@BHY=8ce4HCSD:/e?@+Uf7U:=RP@QV4+eFZUGVI0-+#B.cdU1c5:GY?73]=)1+bW
aO)78ePdJ?MdT=?F3EINe,0#[_,\-1?.]K1RdF\6+RCdJKVN-5NI[0PET&<R-+TX
)^(CYS,bB1P+#BQadCeee2S(E_14&U^fQe3D#^N[3E+/CQ#&IgXX&aefS3+T/)WH
CV_7X\FB3A4U^S6B/S6^K27cFN2Fce+>_.S:9P\Q\0A[UWQbP/,N_?9^S0Nf#04[
f(XK&OQ^OPQe/9&C7(C76_W?\/A=#^7[fRE1GNP&N@C2SgcOQ/>13>5Ma=UVD&UD
TR,E8354afMQa@54LPQY+)4&E<B-E--.(JCgQa32:/OG3V/7EA67HA,LdSZMXZ>Q
Z=?_#EK1N0aO^Vf_.]66@\)#:d5)S0.4#0?;Q6/Xaa)D#IDE^_2Z[#Z76Sd&&-HG
:^e5N@gSB9GN_c82[P#JF/BB2L9EBK1b2>.aN6[ZKXS9MdF@\E^6J)+Y4I(NPad+
4[NO4#__RE7C92^-]&<\/M5(I)aIeE9<XV4g+?GDfSSD\R[OIJO)TSL;B>,fef;,
fF>5&A4J96d0d=ZPeN:c8,/MQ<IX9CJZ/&B,QW]AQ0X8MX9J&B@.[cc6:;M.S>5>
+^+),Yd/)e0O6X3_eMdSBGLTG#HB11ea&bX-#C(f98C2C4VZdRPN/FC<F/bRF-<6
ZG_R^5+>\[7JFBa4IOLRR7X[(]VAPZ(:0ebU(@RZK_&MDA<T83GINAZ^H_YIC2.X
@@J@-HXFQ[W1JR/)QE6S^F?)&&>g/62HV80W]O^2OJK<;?7YJV3U?85d>Jba_]\T
8NgD.OBS6c?T&Z-FLd[][[8SbD2GY^2Zd_SgCD\H;d+0SF6W</AW78S^OWC>gVRV
d2?SeZ1b/gR?6fCdLZeeRB0A<EbQQ879f-gfE4Qd8EGHA-Mc2K=Lgc7=fb6_f_47
75K?,HQ=0XJOK4G(=S?(R2Wc=gT1J?Ne)D.bXK@UA7SFL9d;bH[M^cQ1]BCIO(H6
,d(?f1X#+eCSO^/4O;X4cd)VdaJE.g6.OC5I-S)T^XKH5edggI+5MP6JcM=Y-#9V
3-gBMFZK;b;IF\V:=?=G-H)]W2W<@/X3c86VdAC_A4U[MOT9GHP6R-?UYWZDMe\2
Sg/Zf0U+2ZX^EV[F=&H#)D(RK8\IcN#F5/K^N:a0G<6Jb?\MgGHaRG1I]Gdg9VJI
>R+,19-f:&/+4aX8a>)];Q(8^@f,D@YNF,X\L3aSTG>/a:=:ILM@<N76b8<1R=>V
.N_9CeUU^(FZ0=<5F&,=aW+C?LEG(?(c-HCE^<23Z+?b=f6dK4:H)K[SL0BM9=#F
7^?J[#eQZ:8;7PG_(8)cCBH5F[^UD@Nb5,T0D:HQ38353USFbNVOaQ^[0HN3JdG0
c#Ff8Y<WcLJ8EX)_eX_3<3M3#fNJ(I_a7OPS<]WW6.fF6I&geE/?:#P:>VYPIbEG
#FWPg_\=6a4Y[-Pe]b_5+\=\\3SAG(LH1A8_#W.@Q_ELOHUYGWdSJMf7@X<K\f@]
(^?G:2HJcX..#5WbIbHCd:WYR(]<(EW?^KWQ\8b<&e,5+bN+_(gH&=bYZI1Q87V6
CG8J8ESW^Y0/65UPH6TG,+6BRHXb#>E9A<[/=];=DUSfPT#\4^&_^a)?>7K0_E<]
(2NETJ0:=\W673GN6?::W7YU7F)EJ2;^TSW8)@[Jd?cL2_YI&c3dDM#.b#4FcRT.
)-ZaZC+TLUeI/8H/=FJ^ZS_F,KPEI<VKfBU:]2]0@CN_#L&_ZaW.J78>Z;aE:8(A
KUL2K@0A.B.[6<Q@^)S^ZEO0^Xc>841d@H@-Q47,1P@Ga]Ta7\cBQ>C.NUN?<4Uc
F3AN_BU;d50KUH;E-Z#<IHG[D;ZB>/E;^]1(LQ04B7gb[XEO7\P89OS-RACIW>G:
A0CZ^P,@e5RGab\1_#V,8_@5V6?dfJ^cgW=eEM/W+BVUFOCE1IHM:5=g=;\7>&.#
O_NT,,^b<==QY.][@L&LGeN7[T[JN9JY/UK1XX@\FLV)/1-LO-&+)1N#V.R1XEN1
,.^#F9bI5])?B01IcE3@gE1JEOGCd48;:HbgUf#c0/F8X7M?-W+0#b/cCR#W=M.N
&<WTLQ.7JO;FI;fAX;5g+<3M)]<G(fCC75FM)3M5R(P0Fc3^23PWZNE<D2<^B^;:
^O_QT<aJLeORE#effS[HYY8?:afVb4NDI,a6;3A+3>GV?c(E@_5D^+LPTYN?PGQB
/A7T1V6HE#f.b5VYR)B9F7CTbIG=HZ=-F_UJRDgg15+59/ae/]IY\gb#AMF-KdX,
d7OUI#e5\CT#?Ee#7HOZT,.gO<[F2YaD7XbYE:a4bKF-@?.8)86J)@gIbU-V_\D?
+;>&0X10Bg]G:g0QV[C+];bB/T1.S@:6?DV],,(KQ,73M@_KV5^PJ(g^R+<(P0dW
M;?g+aJ/1KS)7ICXO0QB_@Ue?@>gW\O^N&X4W5<Sa_,_CQ@),:,4W]PRgV;>]c+D
4JQXJ,8I:L-_&10FdF@,cMIIMOTb5E((7@Q\5I.R0GGDV1(#g7\1\4-:T+.g^=//
\#S0b6I_KROM++b[-LIQE2]UgI_#-UQE5>8,AK)<^ZZ9g[,(bHca325A2M4D^C@b
<\f3PMQN.SL/9IZUB6(.PSXPK38HS.X3f->J\f\9N5OI7=-6cZBgdT+212EGP]0Y
Td4[BI[\Y?D@ege\A&>YdFbc-\6/6eUUF];(2/:]-LRC2&_IR3/JABf8a)f>.6Y<
dLI6HS^+U)7&Eg\V8B[:T(=@&TMY4c<+#.U+V5MD^848f,<L;N8;8(\X5+X-dAYX
#)dF_LI89XbF0K8BD)e2,KXWGOK&]O#HbKUe?7L1=FR7Y@H3a#=J,?6P->@4ZIPN
Y)Y&RVSe8>TM:[0;Y1H6_NR3)/2eM&@#?[,E7]TBd54c1/((LV>ZBJ=1V&=1U]eM
3PO)4eJVYbJ1?W@[eCcCPgTa>S296GO<NT2LcEN)1G^#B24dV@O<+MQfF)OaU]g2
XWdH[^K@d(/;9\Vg#A0CSHJ3H&OF/ZAX:8>IAYG,3@AQ9IS7&J)0d8&8DES>?]/R
f2@VDdLd;9Bb5fTfg_0(Y)8@8O:8FJ9#QIf/e9B&X>ZfTT\C(3b19H@:1SOG[IK4
-)UX@M^AfRO[Z=9OQK8Ug5L&T34GS=QF[+7Pd6(e5,MSS2b9<T7VeP06@K6HC^bH
^D;??+2J6KRPUV\UZ\NJS5@bK),OI^&eRT9NSIcWQQP8T??F(JD/TdA@UM5g-D@L
_^Q@BNLOL#PeKSNE/Oa\[ZR&fRBc2Qd8ZEgNf3HH5>Q-Sc0SB+[9181BN1U7R0^I
U3d[<Z+;MJ))1?4LF[bFNVe5QGBZO(,&[b&d6Sg>8N7J@W#W\&Q4OZ9c^65bF6Ag
Q<POa+UQ/FOKZ+[L-b&gICGJ[I,PZXJES^-2O)/N-fU0RRgS<LKfSN-A,?,P:):M
PB-8C<b>e7?()C31.:_,PCM81-9d1SGN_HOaD)M<aQ]<5dWd)2g3J[;>,B(@Z&?.
-&,cOAK-fc\L,^b7WKP^d#Z8ef5#1&aFR)\b)dS#V1:FRTQ:+Naa0H_]XJGSAU.K
:WeR1fdIX^9T=)V?He1<+KD\&-[VFdLH>6d)925Ped:^C>2<(Xa:>8380[G27AM)
_,RC^47(12H&^/ZIE<9c=E-=+=53cV)B4[b-:-(H8LZ+_S0e.9FWC04YdG4^#>OY
TbL3OHDGPRfYTO6dgGS?64=E]UBA8_RFdD>JHOa:ZS?X>P:H+2DM3O97C-SKGdZ.
MU@1C39@L3dEe@6VTD6<N4C@FW13L8=TYb@gXPUAB2\U^RFZd8+T&5RgJ,RNHeOO
C6BWV1QCe,GG)NX6I30FSP\#)D991L<c)S>&d)(Y,=aLfg,)GZ]&J(@O7NZc.+88
SUTI^/RIV-WMGHH\a;49.6c2_0g-g.RN=4HERbSJJ&DOgL#3a/FH^OBSG>bLGf[\
149FQ2DK=cFP-2^2D;HW>I<6PbdK.Q9V9T44P+Y@><c93?I<IM>0c+L,YU71[A.g
fa(O>dW1F]GNO;NG>89E6LcKS9R.[O?HVbR&Ha_^Cc,O,9Y=NPCVQe..<:.5&DJS
LHTZ#2a(><7/2&D]G_/4^3\I/,f<;_H/3D)FB<+2bI2;[UKQGELf6_VO..a&XL@3
-V^2)^U)eaCL(\O6PL?(J/[eVJ(-,^J17Y/78W5L^K\S3EB0H#+S>1BA8W.,O\3C
#g>SG;DDd#M1/>3ad)K(6?1971G-)#F,D9HWa)[QF348Ib@WTLe^<d1>RP-PL;-M
-]178d6\;,ef--B9-<3d/&>>5^T<=LbNNJb1#V3EWgeU2P&gS]c4HRNFSgJB+MZa
-R9M(P@1F/7VT-XdDcFHJ^.d=K._TJ#gbdLc5\\QR[N+_YaX+GB:XZ5Q4G;X^PC[
MZGb+:aAeI#()P\(E71L67QaC>&ZVPU5TP2N<:J1<^&/#,Y;f;SIc_<;3((bdWJV
NV;AII@6&N1U=IDQ6#GXX9ee[WA6/UYcM:d;_QC?0?S.B;J)2F,?13?M,ZMC>(Ka
[.O<4:6-9/=XDXXHOG?FQL81c)0&U^I+5.^\PbT)>/_\b-OQ,7QE/&RYc\I4R_RR
[&EI^d2P.f+e]INBCU@C_0b2dD8Z0&+a_HET:2?=8-Df32bGK40_9Y-/T-X[<.I5
Hf5KaGEHWd9@N:LAb.)d@P?[#\8X(d_,G0-O/Q-gf4&L5T+9eY^4GYE]#fVdIf1F
21;ZcL0@_#_UbK<H]fB<#&A8ZTfeQ7[L4W[/V]>RQC(g@9]+f:Tc@,P\FDS2FD+X
JY4gd(++L[9=JG05#ag\T^]1\+R]2Q(:ZBQD1YYC,^R)aGOM?;3cc=J4JJ2:8A1/
e]Y,<>8fW&Q\OP)-7O03ObcEGA75O]7.H3^:MCH)1-Qg/P\b.VJ6:f((3d5SA45O
@5C.>]CK+<>^&]\e/Q]-gXH05.8E4+(T7<O]&M\;^X=8QI13[EP2+)2/^VXH0dL>
L3#L[10W9@^)NTEGH+/@MTg-,&L24Z>)Q54FF5b&B_KW+EM6&,\f=(aMSgf.IWNT
JVfDE7M=gO<8IB<NSU^YeEU<?#]bQ=XY)MHQ-@HL/7#aV::VL(edaV.OT;1]/6g_
Ff_f@LbZ0EJa+SS2H&TRgUHNYNBIQ1REI#5N04(BW]4Ng4eL4T0T56<DgV]\f]WV
5ERX+.J94Y6LM?\#<I6Z_+<^6,fCG_[81gQf8dIPJV&9cgfTUS^NSeH;<<A@IHC;
1N&F:&d9TXV>Q903TKPdIN2FZ3]L,.QZ[B<Ndc.;:@b1bL&Wf1f<_.]#K30_L6T0
fQb5e=+,BXGg[K=V(?83:1X507&(f<XJ;I_Sced>@dc_JOIaDEO#]Y2@g\G;:e)6
4U0;1OH[W&(MJf&1NJFU2cb)MEDIAgcYDCIaU?7aZ4Y2:8+<J/2+/D[T.:72Dffd
1O5?5:cCRe:>(ecd<7>+J;K0:K8151e8U[[6dF1<PP_M\D<ZEY5CC-FPaT<#O(&\
8ZKX?2(JNfJDO9OAJ\WSCU(_JJFG.OD:&Qg6ERF20Z06K/8TW@4aRI3Z-Q;gP?cN
H3_)DPg-gRDJQ1&LT973G8U7[-a6#R&OHZ@@XQ\_J7HN-gc2F-TbggJ?HX6N)PMd
PHF4g9)dRF.,af#ef?F[d(Z>:=&cS;U&_L\Fa4K)=]dYOLL/6A9X6HOc-AL/#/\(
W9bb\KHL+6S,e7<bY[)Aa(D]96G+O5=<e>-+>AP5#4,_g18Qb=&0-KYf6#?@OD^f
0W\@F&[KKc0X?52fHPMT][eGKae[7,Z8d@GbP:T8_&J?WgdaI6<G>:O]M999Z66Z
B?b>S,?@a<aXP=JaI0]TP83Ua0>[0?<Oa178GgOC6AeQ9a@+@=XDNL(-VMC[eBc\
gF5c\?_I<]bFSA1M>0#E315^,_F2GT6_Bb,MJ54g6+fM-GcJ35JYC?+PTVU[.W6&
Gd[@F4c&V/L+G-;[WBH>A#O[AJ.We9^MW)VPcb2&ANbZAPO@YG]+E@40a.>@6fN2
,([VU7OD0V7DUWX#>4KCeYaRP=HA<EPaT/&17M;M6(MPI-22B\Q9>08]aC.VL+^B
-7eTR#SL)UAE;c)49C[.W@3[Y+^f6C>W2.LT?JI_Ng<R)(Z/OcZA]c1<a(#Vf_c(
R@EQA1RH)6#OZ<DeJN/-a5FZ5Z?R^4PK,F\34fB[Q9\P8EZ.Fac-EO-RCO[NOQSV
I-8/&/TI;>e@dJSC;O93g:#RG0WD[OVNCd2C-NL[8L4H;7.ITeb[eR7<]2G\K:Jf
5H(TNVI58,P9JSUdZgB7c0.TEK=6R<AI.VAH#TdBH..1X4_aPC4DB3R/&R\)D-4&
^)&Y9(W?.X(PFQW>LR7?:bXcCcVc6D8ZUR>K4-V<A&J7f(ag8Q;+DYO]?QG5-IP&
Ee69cOfM/F+/][?E+a\EN-#ZLBHe&A402/=@0cH3@(TN#IF,9)beRC:)S[);R6K4
+SScLD;(CgNLMc+-5Tc.IL3?MP\.A0f=1WN6Ec8SZ\Fa7EM\F0fH@,F07BGPcB3_
eAOK0[:S88;=edc(E5P1D)NaO+baM6fXX]a,K0V[&T4WTg0@>21c7Xc.gV]S-Kd>
Z3SUE@G6Gd5b&^DMA:O07K/8MUM>PFfV_)<_8\H^W+81@Ka798YNeJbOW4#YL2VI
>D6]U15MPR>9V,<7<VA\7M.Z),32T@:1ZIcQAbHXg_Q6fcVX3P[Ua_URa8RID^GU
J(:/CB7YV];QPK7+&F8]g&^L9HO\>eG)>H)G(F8=LH:Hb,V7YRN<eAMUWJ2F[9CI
_IXfWQ;\#f;68B^\_QP,<BK(_A,Q/E3@Q@A<2AWEa]G;1ebb\b+_gV<5XVT:7FKU
bIdLE8MLK-X4120KBRZb(a9bdT<8SLI)TcSV#[d;/DcM66cCI^#P0e0PWeP1OVSW
<]UaNIf5FP\fT=F=WNc0eUOMC9C<:&BcK-B\Hg:Yc7[.fQ17B[R?<L5JdJ/UH4c7
OfW=S3Gg?L1fRc-4Z#5PJ4K)BcW@<>8c-YdC#>V7?U-_F8+_QGB>OWG7gf-/7#f-
N?1-ff^C+,J-&-a#&#7B,/58R]&9:\6D[Ig_J44FOWH\KZIJc[ZR43.+]:Qg&^VH
TXYB?<KgJ@=.DM&d,.5TVg=BXKO\fSYgT(=9\BMO[<W8?7PRW)NEOU\R)6GK_9<.
GVZLRd]9OF/G7;FL<]dUMJU6.2[6=aG>Y_0L,6=A0Cc&g2F7VHS3:20AaPN=6>T,
AX;<#e4Je3Y4f5JCS4)da=;,TTQQH]d<SVX6c@d^?P2_BB,PJNP[&K6d:)7_Gd0U
:RNdWc?UCHKG/1L;ePVXNga,E3)P@6M=#9V.c3a6eYYJCZYd7>SX_)eVZKJGAbZe
S#^BY>1-\bZV2b=\4c^Se[G<bLETReVJVT.D;_T^UBOK-c=X#GB>O)O@2+?KQ62>
IRgRN.CYP0WJK[TYN:d(gf8\Pc\)<8[;U;@6VbW?H.QLOF+F9Ua=6WgT8\Sb/Pb7
7^3:IBfXC+E,8N+1cCJN75[\P/4dJb#+E<N?EGP=(]g[G&(=d_35AGfe-eF->4fg
Od+_R5c7Yb,J6[_Q]2+BH#0IUTQD3#bC0OS(3BC1+#O]UZ4CA@QPKfAN6cd9H+#6
DBa4-B#FN3B_f6U<H);de20S<2PM=U0,UEXZH/H&9N/BS80/<@.6TI7>cNZaD@QH
2E,,=?[83\CRR,+T]>-N3fQ>_;f&4@8^]68UI?VPc+d+#\@DL]?5U\QF4B,EXbg>
TE4X6Q-MU[Y7KK,[\6YPM]:F/8SA8CK\6N[BWa;g-7f-FFEbCJ>:>@X5f,WCQGB;
3@5EWg28WP.fa&L0\4PD-+<g[YO6-A7OY5@229T:Gb.]JU-EL9UIE;Eg]/ZQI=6g
2/G]]U)Y9-C#ZPTY^/R@@=Q\@&ZI:)AeBH-4d4FBLJ\:O2Pg9V1e6d>1(LUPE.[?
EeL8ZYe<<:6dVeJL.N^?JV@C]ESC2&07MW.)YPKUcAX^Icb58055aC6?V#?Rd=-N
G,3+M^B7#Fddb&SgQ3QB@2KL[EM0P)4V:Z1I)SIFODdH;JHD0I[3\\4#5cg59/L@
5-20&OQPG[_P.G=6[3B=f>,#/EOf:7XKg81B4AD8L58Lf.#Uc-g88e;gEU9)#GX4
A17.C1MEeM=YWB,[G3X862UbcZ92e?SI8V.M-?g8e_3L5\T/?eK\D[^@=]37b#0A
a2:6IVbCZYOVN@@@6(/CJDQ51c68^g7.,+E0@]#bdZNZ4^cWfJXU:^E63JD16:)Q
QL^AQ6B=6DGPIc>FNX^<M8b=FKIG/]>gVAS.2[(+O:J@(_40[_^^51EE,YJL6E65
1&.#8=8M^)Nd38T,:N+=#>DZbL&Ef?(WPg4:Z[g;QO&384Xf4bYCT#O2EE8#bWDO
R=VL.O_8>Vd,0\JR:Y#L5&Z30;E(]-RY^HYH37WB8aQa?1@P+XcP?ab&5)[5VBLW
L6&01,]g8(^<&T3DIA>/2:38:Yd^P/aV.0@5cXc8PQbZ&8>S75?QEYDO21Pb/YM@
_5^Y7><4DXVVK3[Fg[3T5(HO;BW#_=C-(1+U6VE8,GJK44KU.D]N2dH1@W:(Hf9M
AQI++>@f?/^.68T22[31U7cgF^X:PUF@:Ra@8eY63HD5=^LSRD77:X;KHEec,CS;
;f,)Ze<FSWa58[H.V#;dABdN78PKMNC6efUW^-@Zg--9S:J^\bBcdE9OK^aP_XT,
,e/=ID1A+\6^ESJ;T@>YSPP,MUZO@&G&UE<Bc?V/:df+5,QZ2d3_PdVJ41:C7gU4
\I6=V7Edc2VXH>QH).2>N8A,I1E4IcOJ6AI1\((BVJ3G?&)LWaU@S=+L#f[-bda<
WF7^1Dg[-f>WLR/SLQV:GC=P#Za_T3X8EcK5R21#&L?B+N-(1:->4/2HVY;WdL@;
KNPgVJ#fCa_fN->bSRK<V,N2CKXDQN?^T.Jb\+TRZ(XWL&>.F:5WLR;D/_+=4]2&
E(>A,4)R_;?WMBfP>@#(f4:QU\]>]),):>>58<c+<LAY5+SIaA;TEbEf:fT]A,@1
LR0\J+7fJ=6.CR09-DMEBVV;AUZ_]=_8GFM_L=W411]GD3(7VOL6<WTD&)<<1;#c
@\bC@I6)0KBV8=D]YC?R,ZO4Q)Z>>f2C>KBaSOQX6&H4TY6@(2+2N,cQL<P5B]9I
T@ZDc.Y4F:HSZb_>AZ^Y:fY]3e0@X8CZLC_/:\&;4T37,f@PA&NKY2=BFb4)7?)Y
#XSHGeceg</ZgdO339C:VAaW(cV33N#N&aO)&-\gA7R0g(/0@d73H.XG/#NI>@X;
<_#]K5g/106GZ5\>?+,#fC?b=L\T.25RJ6VQ4d9MN?M/W821^<I=Q(a6P;[?OF9.
DKN?ET;Fg@F)D4)UQ++,]@S3=#JES.=_J45R3)DRRNf1&:L).NX:)bP0<d(dPC.8
#;W1CJ@FbH(-Y;5;O?-;&NTQ)4T8\W^a25^R?<VI]7:L[]\1M@@>[HG2dTG#T/IM
cfM8V>@M#&/H:99Yc>g3fFRXYG)@>L?eHJ:.X9]#/4Y&M]KJ/VbX5IN\#>?f6UHG
LV>_8_TGCQ-J#Aa<O#4ER8c\CVC@(AE^.FOVKK-?IH8\gEJ]8-<9MYIB<6ZH?L#b
TMdF&gPR1Yg8,)Lga9Z-<Q&KIc=ee<DNL-Q5MSUBg1,R2FMUJ0^N[)O:#\HDZ?SD
.F+8X0L#TgMTaG@@G8O/)6<;(4R=,08_eaa4I]DERcG+<<=+-3UT<U?aJ1g5g9O\
26eP(.L77(15,KI[21/IXX?BH)+fU=KOW.,)3G-2)G2LZgL2W6d7<_Sa>eaM_4+R
^93:.?ZaO_IWe)Oae+8f3)EZgB]?_^BU?CCJGT>DEC(?NdTB#f4JfaOZB@@V^V[)
d321UB6IcD</##7I=gaY<>g\W?g/;K9[SF(E#eBY>A^CE5Cg&7=98)P@7#3QGHHU
2OEUTLYaaXG[1Da2O)f\dZJGI4Agcd5#UB4IMSdXIdI5C.48\C5?UYDI=/:Q54b1
LQ1aLg?K[G/&SC48.g@0_K]\(YXN[\I,STF-DZ,VP,a[)X-GeYL-I.a.<FD+LZDC
DFA](2RZT^9BU++bNLAK,XMY6N<90ZOGRY&cb25&8.?<96ce/7Nd#GN&,8KgI)G<
WYP\AP\7E^6K(5BVbfbN-.cQCd0He5OBdPB<HS>HG1(30T>+C/(NCOT_V[7F-S;A
c:P^:-QQ1aQT90FTXbP>H.G&X@dO&C\_5KQ&H6=_+#@SE)aF?4SPUNYD;fB5J2?0
UdV\82UR+C&Y;^=CRFa.^7)c1Yc#CeH_#=0_I;PE(Ea2NM.ffXEBZXKTTfA0=Z7&
BWSXaEagVA_B(Pd^LC4P+K/1#><T/d_6>:>U[K5Mc+U\^MYV\.\:KVKM#(:;3g3b
O/5>6(W&>aY[AAQ74/-&b0M-;8P;:/E2-<]TQ=HF0S]a=gX[],(aFgV<ceMLLf9N
(\-7f.e:JJCO,DNL_G1cWL3O4&BNJ46H(M8J3YD(fS)<Y=e[3EDG#(N?NLb+J8N8
MTf-3d2X:_7d&e>S<=YRg>gP[RI)0):47Z@>^;eC/aR^<FZ^HVBFB8/W95H4SRbC
/5<VOF]-DP18[@O7I_>JG&81-.<aWC:Q#>fD&WR6WaRCCJ9IX-;,V&[g&6;H0C)C
N#3XDcbA8Q=bFH[949eEd2L-Q)g<=@g#4)7+6^bGCOP?^)>;,@HgVK76F0U^XH[F
NA-P#=G]U_9@/Y]fLJ8//;cF==S4aZ4Q4GS[=L4GW@4B]Y4U\0(Z46?g\_fO>Ed^
Z,OfFUSMgb&KUd@C]GIVcT8XdQ@e86M;_DY(V>f2L>?8>--_[?P.>#LM=UA_<(-E
Q95EDG[T22V/+S#+d?.#]/SHM8)B61SG2f\^Y<RbCG\Y>6gG<aC;8[Z@8@=TG;+P
DMWP7fK<.V98;aeb&:KcA6S)592)cD^=ECdSfa+NX7#J;Y4PDD=3CQYa#\1bW?_R
(R>)2-44&1,:\Fg8f=I4HW4YM-QbK>,X3;)b0;+&S03=DW9:M9.Y:\R5TaFg-.MU
O?f]_febfCXSHefLWZ#R28f5#,:NA6E(NY2GCHEU7P3&_>W_,?WPTaK,JaIe:X,D
EOK/EHYLODC]0H4@B0UFNZgU,1<U@/^(T+>EB)&)g2B3dVJ4+c&g(5;Cb\23<2gX
Y@eNIaH.)RRA(:LfB9da=^NW;._.ZX3LO:LKF@]2([Q#<9Va-T8b(0fgBMH/,bCU
Aa@HDZG]M-^#&LH@;MEC=1[GK1806Z\]9VZT]C[IM&=^b76=HDG^ZV\->IQ]d:I:
+>.2BWX\MRXDI(W22(Be9KFa:D6)[=N5NCO29FE>P.Y[_KeCA)H_Y?<g&^XH(d[D
B[Bc0Q#UJ<S:-?Oa6)bEgI[UP(PL51PD-KPD3]JUGZY1))e54TfC-)9FMbSgGV^R
Lb,6UDEZOXb-E(DB.@4:EP)^ab[O&^IC7e]A1,F,>2^@.U_/.^DFXD.64J=;Wf3U
MaQ@=SW@DLd?TcU-.62g[b3T=c#]DJfDd\fg^9B7L>+9_+F\(#R#&A@G]YV;V,.2
cCGTb@MffQ6fd.NJ/0E4__7D3-M;7Ob2G-H1eB\PSdW-,a&]bfJ/FP05##aba-Ba
OT,KSC:,S?>_ZUG#6]?a=AR,V7RYFZH7\JQI33JX208Uc&ZH.<S(J_cB:>F-VFQF
HfcecW1(8],A7MYJ>YWCS?^C,28#cLec]4B+?W7?dN/aWYJ1TKAXURQM0f=Z>L[2
5aL)BH.gI03E9>EQY_0YP?a=LI[)H7=[OAI^L=VCd5g=0&eRA/4H[e)TJ<HO\L]L
5&?dKI9[&@[F/7^+(L+ZTF1N;,RZ^KGBP0,UGbG=D>]6)O9I-.c9Eb[2PZW:L7;P
,2\=#MFLD60/S7XF+ITJ/V,#RXKZ&6dC1GccKL;@CD_+_@)/M^GG]F;^<7BNdT40
G0+35]ORN7)E4RaI#g1XXZ0<537+__&12K#J,-@;5L0;D5<_]2RLVL0/)^]QQ[E,
8bAI[G4B,7b9,.P&(&Sg?WYUU<[+QRg6RO,<2TK9TfLPKVYZ,ae4ELGD:7VZ;7RO
[.N,FbGQ2;UNK/0JdQY-;H;/1,J:)GO<:/CWg\7\f+ZZ#(E(EbM:d=^EKKPUNJHI
^&4V6M(;_M91:3/,JS6FX#e.-:Tc2#@Y&XW=bMAaV::NbC:CC/e+(a_CUD44Cg\&
P[S^fO.f<?2Z_<;,5fgDc=9OVO>NAJT/aE561ZVaBI9,=PW:3[EZ4+>>NeE+fR.O
f&8L^[,bVL-?#c_@)7SHcJ2PC&PJccg3(YFV).V+QYG@H&1_=IGZ-H;-M6^0,^??
_8&eM-W0/N/1Q605=C0RA>g(<-54X/>/7W8AN[0M<-/KVa,b>1(D]2Q7@d:0L?Q/
a=9<7[1P?X3gL#8Y=ag>O2cM2:(Y/:VL9XMFDS<X5W>8+;X-UI+(;BRO[9adbUgV
,YSfF8Ab^U+[,8W87?ZK\a6#T&WA+V?_/184b_M2]06@KfTYb<VVIC8a.f)P?CM\
7-6(Xf[12\6]AdZKV2XSK69()\[4-VXaP>##E<@#4<3bL_KFJ)Z60dT6N)DWdfaM
T,&(4c.S).I>;D0KaX]fO;d=[(IS)c9D..>dZ,;COHMF9B;6P[_/g<FA+;(010AO
_[<3QH6?]_>R)=8W55E0_BYaeG<=W1#G:N/V5g5L?/(SGE?3-8&P6gFG.I9ODO/O
cb-a5[.CWLbJQLMgH&_gaOcP-H3=??>BP?1J]S)EeSW:f(gJ#R=e.6L,ZSWS9Qe>
>ee@-?_HIcX76WEa#,cUDLB9U4/]O(98:D&3&88YOD,OFBL4I,NcR.2eZKbA44gG
W&3QB3abbfQF_c&:&bb1D<;f.UGB(=74d<HSFeJB3Q4T]9>1LdU;/L4OMRZ<J/4V
.<AJRE/F<M45+c/D>MZP=@\N#N#Mb?P?6<D_ALc(56RW_1EUcgM1G>8ZA]e@[e]L
8Ma)B056.d>-LL-O[>JU63f^S5VE)Q4A5P@]Kg12FT^BI.?UV[+)K/8\ZSL8gY,Q
G_]64Qce4EP5&8_R):,9?LHY/7GF=X@,[IeS2_6H#LV^75:4QHJAEC>WPdECS:Nd
MZ35:RW1)ZV6+HIA\H)/b\Ve2dfdKU#SDH>/S0/?E9&;E?N;RZ99cAcID,9UQ>bW
F<f7#1K&f3#7NFY7W3LG7Me;P?=9,RU?U_Y6Y<RD3G6P8]S6\SSX>74=G=M>S)5D
a6/6WIV2,dIJe58]CUNegbUXe\@@DB[ZS++Y[XU_?c,F]]abT>^TU+RU5+2E.(OF
d<JGeXO3.-XbBIT):J\Y&^eLZc9b:9DH^(\1((1[\c3C^>1[bVMJ.H[:QI4;XU_[
PY]JJ^R6d^f?>U0@:Vd6ace5Xe#FE63,>8f^19<?_,MLDFf&g5GCJ2F?PfL.2<+I
L[E@.QH7Z39Ag7TR3S3O^QGW_EIL^8TH<N7NQ:W\:7-N/TGdKPY)I]VU;HOSDF91
Ebg&\;_[1N3,&-_G-FbYNUJOa#HD,KXfgB5dKRa:^-=7S3^Q&(W:T02=+,HY+S@:
A@J&\d8dVfAE),2N]]KK>6=5\)9gBC20c#J7F<AB>MTI:RQ(<_NObXDON]ZP#EEb
7^=@c:-30bVVVO.YE+dEAeeKSI2VQgJ3/\VW&5+MUM)^::cVeH[Z4^((>8?0b1XL
V-d7WDbbX2)-Q=(?SNB>[.E5U2[,PS#Y^dDPc_/;58g8)b+c&DN:(f4H5Yb4faM5
&AO9A0BQ6N+?DU&F(&@S;J^06-:f_\9WB^,eQ(.fg:3>B+]++YQQ_2/&:T>+91;b
V)RUMf<ED:6:QDU7XIJ7,?D?V&<.,W#L,8Ob69:Sb\FE:?ZB.SdK5HJAE;GOd19G
TNYLI>\6Y&)eTbOM5dFN\b3?9H/I:gc3.4V>aK(2HD\Hg/7c&+9PUbQB/ETKd1G-
&cb1N+):31K^,VaW;UZO-<&1&Q52F\FG^;YYb]NDDV^g]0X27g^X>7fa95Y[<dZ)
?A_-EH9aQI->QVRL-EN7)@_U\/FEf/(FU,/77)NbJ@[IUJeI_?.0PF7<cd12I]8a
2@cf=RfXMW4^(Je63XgE(#?+d)PgDBfYdeKOdF_AfT,:SP.3@QN;D@RF\+LEW\Jf
\Gg]AM>68(>+3@8^DI0-e]e#(IH]d[IT[ADA#fMRXM?bUDJ-SE>&0:(N9;CB_N+&
.CDf58PDA?]1.19U@(F?VDf@F^^5O4K3\Z8F6&6GK:E3L=EBLbIS-;cN457F[433
TB]04A]J9d,UKLTK0L-If@TTU-#1:DVb48IFN.X0835O91]Ja6D80La=^IfX8T6N
04Y2<GOE7>d.-4BUd2=GH5.[dZQ3[AG_M31P>6V=P.2Q;HCAS1^]Ig-)])Q2:Z>O
SNc75^1SGWN5VBJP[8Ne&N<DJ3^318R#7PBZRa8J@\==1d,RV@(bK+5WdfBL\/dA
.TS8)c4XE>UUY_I8DY,\ce?TUfYF>9I9=3PFLeM1T,<M(=LH/HX(87D.A9gIC>[K
#bX/CaH9=5=KO>f5fH?H376JJZ72O[+;=B/8J1>84</EV)\DJd.I&>[WIHEN=7c)
TCC2ZMVGXME7WZDUOMf;1@+bf]VIK0LH+P)US_d\A.(P1C;.J&\E=4FA5;/O()]f
<G)ITX]@(#79EXb=G#1K7BVNR:Re.aEfNMW:.d5),edR&0)Z^Q?Q]27f=JF3LJ(5
b8I[L9Y5O]J^2?8g1+&9:OQVDfTH4WY7;Ae=#,]FTRd9I@JRIa]#\MgQT>8UeI2H
(<a2X4)+QC/dD+V1LbE37N#;XNV/&E]]>^+/-\UM6GQMfT^E^9_7O4WNKGRK]\BD
]L_^TD/KF;\N6cK[YTURIWB+12X]7CXUEYYVBOg2f@_W9Z\G-X/]\:Ea^1:-#Z8,
N0.E19C?4Q]2Ab:_BTb/,VWW?)?,13A5bSB8Lb(35PCQVFNJZ,Kg:L?47AGDJIX/
D[(BL@XM[D,=JW&5L@,b419&(M>8._5;)JGF-:SXd(.?9I1(L.F5-/Z3D&QQT&3(
a\#Jg1+>E:NKD&&&fKMLBY9=fHG?b.HB(f;3Tb(4UDPWV)5W47I;UGeB+0RKWA[f
[4V0J&^#][CUX;=K\@.e+(Q[X+a+BWL&P8f9Kd;c<IM9X?7bP8B<]gXO\HUV0EA.
DPd=8?3(>ce0<[:ETD6)ab0RLUT.ZKV9M#6g.3EDEPT#S33[;5J3JD>;C)d7W:#\
d\:9A=+bG3LVGEe/?HT0YYd;0;3)=3Sd_TdP6Jbbd6ZZ+[1FcM0-Vg2/6:J,,NK6
PD&=U&5PeU>WL^=cK=&M:8T/HbH79=68;b:^d50O8PBgEc#Q?]&JXVNYXI:/G-X@
EG,1_JTCa_Of.D<.;VO3;V,E;>1/,71EJKQE<\bFIX3+XPKR#d49#<e]P[4^0I]S
B[H9[P1AbA9-P5:b_95CXK4&^TZa#7Y<eD91@gBN;+[2^W[[4S(ZHb9A7F0=-46F
=N:.;b1&GF0606e.[U;7A)MTRP[Y[M=]:32_c2Q)^IDPJLG3aDgWdT0<SMgW^6e+
P08+g5QA^(c+O+a-a^GJVDV=8X6FVQ)._C>VEZZfaVGB([6OSM5.\0Tb,3#)]<8K
(,V1H89_Q[#KNFO.3e\+,?=VMddXY7c&MTA0+YRYeK,(AgU+0Q83X7-C&Q+>F?WE
_+D_8<6Hg,U78XS,#W33XY\QJb0d^.&@OX_UIC\AT=954U(J93X6d.6,6;D_5GB\
8F(Y>8+d8IT/?@4GGV-P6^@5&eM_+.Of+]4;.ON\NK;ZHN,1KB026/8,>VPKQSRZ
?[I/4J[c-1QCBdD5L]^JOZEUU8cJMQ4=26I8I16)23P#KL;K>2_AXUTd^W_FJY+S
\GW\d=XU8+L?9UY-Q0MeZF/F/_[5,7+bSY0USO3J@^64d>\6X&Nc-PU9+6(^A_OK
S^72_@6@S&2(C[gB:bUB:+DDU>Z,8dJ<=f9F4@>GQXPbIdBIFVJA7<=EP_P)ZVf>
0.VX[1\FD+\^#W5eNSW=0BWAPEaCFGZ\3gbWWYAVMJbcS6GgaY\J2We<Rd1QM/Rb
SXK1)_2g_)?<>g<YZEe]CdC2-Ed/f6>&_27O]R]9&dB,_&7@UVb9J@//N0-05GfS
Q5>XZcD[d.:@5F8/fg:;fOY_;MQJ--VV8&_Q+5VFBK^aW<OV)S6NE8V3^MLM^Q.0
-U)ZIUg]A#_^5egF8L&.)Y)bS7&\(EIN[P@e,9;BgNgB[05\YH#3V+WB=U,?K)4.
F^:Q>AH[\WD17QJ21E0],T7FYcM[RcebZ)/F:;[1FQ?=.<Z&[60-QEUF,+VTE3(1
:Y9=A.6-#geVG(H@>IG6cKX;2][H9T?bb@0/DS4HaGDT6>A#=S5L+D,HdO7J?[^R
W_T0?]4-F[^c.?+]eJGNY..(BcEeS&CKIaF80#V.(;&NT1Ra3Y<6QA68?W)a/Z]b
b^a>db:I-Ua-)M.gb43e]b((,C9/J,CA6M]SP-bP^eb\?AMYfLD+16&_B,.30S\+
Vg^@(Cg_IIL&VRP747e>/H_8_gf1JQ[)D,ef?NCPebY5T\g)F/8?e8F_Zb8ZE\&I
7OPVcI/6e,5g+gJBQ;dLLY-M^Ge:FUaLI#PRe/MTFBXPSN-dgRYPT)a[N&MIRH6Q
MYd_S(-.W4ZR[?/=?)\DTT=[Sg]1E1b+E\d>.0;&e28STN3fFfff19LQaAg8:Y3A
RId\,3;]1^9[cVAQA>:W3/a\,g0)^1Y;^RZPU65MQ]ZGfZQg-HU;A5,B51@AIWH8
DE4e05[AAN&8R,9gQ+&U\Z.bc4cEbIEf9QFH06HMQD>)_K6_LK0KVQD-a(78M7WS
C#+cRB+WCECVaNe)GAYSG\>_e[[?J;e3^HP0)JV/]_@(NcF>1=KbOPg3@_&cK>L5
aQBSLGJcM)0FRONSZ],1)7Pd=Z+@D)G;RTP.1HEfPfUF>;=5[2(EdWA8#X4Q-RX@
fN-][S?6^3^cB\<K8G_I^M5XPC-[&)\5UQ5;=55=_::2X@^Q@GVQ<N9OJ0G7#G9J
e7SR&ddeY)P0[?NMf.fP5?UK6C^XK__5KS:=LUH_>FfJXb3G>IQRR57A/4SL[3IX
CRb,f\EJOaZSHWc2./@Z5BAPbf9GCf^T^#ZCMgIWf&6\La5,(H<#aLV/HO]J@H]H
If[aTVB(^c^>c&I2AbbeHC:Hg^c/\S>=2G(aP,\f84c.afBL0\d\,6)W8,K^G9&>
O>cDFMHG^66C0b1DK?;R-PO()^Jf=I+=6aGBeG&^SUV<S)Y-\I=aE?8agDVVTG:_
OD4^N_d><gSSaG#J@JC[7G9faAPBGGES;2B)T6eLT\N#Q6Da#KC:WR^4ZM0;P4/3
\5+0(9eFFTfD)DD2^88IdBCK;D<X6EAU,)D[GDVW55(&#VZLf<3cQZ>WE&:c7g^#
]Lg]K^RbQU,;GY@,LM1)@_91IEP^0[L>\)^QI9NQ>C+I\RK8;J<W?W:\2S,>=@>c
<1B(a9f6P^_IU)Lc(Y(1YPB84adF[S3PMX.DU1>/G#Rd4Kb5^=A8A><5W(O1R]Tf
M][#YEZMTRfd&1,L59<d#JOL=E[S]^1^UG:>F;;F?Wge/R1DI4>@N:<>XIC82;K+
B&RO<XdD,G)03@S=]J2cU71H9BEB&YG;/3CN?C+Dd<gY3eG)4&MDag.Q0OQfGL#A
eZF@N2[D)G9A1\VQ.:7\POI?T:B2V\3P[=17,0(f/cE++^(dYLMM(#QGReZfM6cE
RF,bTPcG67;^:R0e=]OI+#6104E5SE,a+^Oe>W;29W-8ZG8c.cJcPFAX5+b<9F6@
\:c:,EL&>_QDQRQ:@?,cQ-)S0e6QgaE96KPSE@U6f9=d[1[^7Y^RZGWAd?[G@14T
FBK.6X_U,e^3Cf2+?Se6X:GQY.&SQ+dSUbWQ[?AcabcC)<fK?GL6-<V-<QBg=W[Y
3<Y)X-5&P^R+@VTU,RL_PCbeN<42aFUD9.?gO@V/;5@J7[bC1W:VBTVS8C,LOIB-
MLEM(--[JeBNBE]QX9F:X<RW5,c#C70\,8C6[X,4;G2)M>7S4)XNXO=<;)&Q[HZS
(Ie#M8P-DP6Ee)CWP:>FW.UD[3=Z[M:7&0<4V<0-]BZGV.<X=SbU,RM12F@4(J1E
RV\SFHK-SGKgbA2XbUH31HD[3YcVS7Y:10L==1=:+KfN<V@O7C:6GVA.ESM@B+JH
;bSIF5e2@5e1f7E@1M)7B<af_ZKc9a/9M_D<[Z_e/D_C(NT4ZUF.#X-[VA_GAM08
?P5KIXA(MB2:d.b+BQ;I+37b2.H@PX??3)eVEEf@:2CINI(F[UT2;ccW/8<G_+-Z
6c8H[MX]e5V+OJ\SJD<BACaf49b<_=O\<&;O#<.^JZ(LO;5&6Lg@L9ZTP/0-?96P
+-\(O)MBE2fa/::.;5Y++]IOf)0?->)2b]dME6E(fW5^-d[JS2T][YA,,Dg(9bQH
8/>>]UbcF/MecBCCD:GbX?#7OUXf?1dFa[T78/#.WaN&=:8CD^FHgSQ,[CNANge+
U3a259Yd]CJ+M1L1R:bDC#6d=8;),WF()gW(#I#\JdFQV6M2A:AT7E#[OAAVC^e8
[[)#,ZgI[gVg\TMaE_4=3V[F)/1MC=?@MLS9:aD@-0aJ3X1IY\M6dcCF+/Y,S7;E
-S,QI#Z6bVSTJN>ZX,?AO4R1M)NgbPGY#F=26[=PBg--&#<RAD>J@^H@W)+4F3;&
3NdeWR:Wf-=+0273d,IHIMfPG.Xd\XdD>^XMD(+bfSF:>N3#D]_=GWN/bI&\[7Z_
2EM5OA2E9/D0CdPTMFZQ3GNbdH3_Z@O<eBB51JXWQ&VL3aX)NeTJF]fP)YE6I>](
e;fT9Fc2UDgUPa#V2HCC7.e/@02F_fHdIY<2JYVKVG#/[Fg\48=(<87-TZ(.YI5B
?EG32\@&AS0>f)gO_=K6C;0fJcb:<6+?gaTaX09UX,_(cg,E+P;6+(UC(Q9g0#RU
GcJd\\6gf887(3c793J,7>BeCdbDFZ3b]G2:D(O2IeBJVcd)Z(R#9(RY28K#(O/4
QI2<#\4YI.0)AC9R;@98?.fL5),E7GYe)G(-[,<WBK/CGf8g]3SQ;G^JXPO]CcX&
BDJJ#ZSVB<D:OVb3[WRE4e^I:MUJdVDU&e-RE@GCe=[YEE9ODa);NRN&Y&,\<fIA
b221\-Q:9G_;S-YXW:S+e<LZ:ESPPM^e+D7[YC;.AT()=]5>1;(e1aJaJQ<;)JEY
)OdQ<-2HTG+X7^bC0RW&)QcM@R&(;X\</<Ra64(d^U<F-+We\8(3Mb0J=PX>L,=I
J-R#eTDXN[:_EY1R7^/S24)b^WNUX7:XY47->9YVESPDdd:<+#8;HCR-IF;0<Ub0
O3=C[UUSRCCNaR9]e-BYfe;9FgB2DW7D4##cAH/Pe(e^Of7:KZ-5Y)GI>8R@R540
..XD;CIVKJe;/ag-\J:T;2A1],\Q_XS,E14F:\42J<S/N@VJc593?SK.W&ISC7](
><?7W@(eHR-UV8ICPGJeTES\./\6-<c0VDLgO##/ENVSgaM6YUfQ(S;)^b(/.^g>
Df)K,(cbZTWe23Gc<G<@gSZU:?R?V_]B-U.Q>5JHN7(@8+(/4.&HXIC^3B#M)[00
c3R.F9GP4+8Ea^VEV@.#6a\,JR_?40G^RH:2EBL+E#83<#2:/4?D>+:9V[NIZFeD
GI5,Wd4&:bIa-H-4)/MJ8De0&G5O6F;OPVH;;KU>+GG/)P@NO[7Q]03FFY0<\-,_
OSDV\>F/VZ6XN3G/WS&FN7&X1aGO2Q;dWW6;X]1Gg+2WQfQH#49\,QW/-^.7J3c.
eXN<4@0)RO)UM&N#G6d1b8P811fSVa=#d#gd8W5SK#(TLNOYb9T<Y=:3a>>#Uf8-
O=UET;Q5O,=;;cdCCCeV?FQE6]ZF4HfgfSg155]#@0ERA[/gPFZA^d/7ae,8/e)+
3N)P:Y><=dg8);gY2eBc@6=?T(eB2V^PXe7)a5F7F@Bf21)(Q:426IKXKCfg#@R+
?,0QHdG)gI]3_&QC0^5P^?N>N)TI/311UL>-N//HWHFY9M9BRe^L]4EW\?g<d\C&
9(3eSaeg:CZ+P2=VLfZC.M4;(JABBL(14O+Y>7/;Z,f8^1H2aT>VQT\U.=bZBFcf
Vg+HegD()JRb7-TS3>G_LQ22(8/6dJB_LH>aU_9Fg3(O:P[ITJ3/E1V+DGfICHNU
ICC?1;1TR1A>=EA3dd6B\XfZ&])c>CVHVA>73@eH5^dcB)^WF_ORF0_#DMI]X8:1
TR&6d8-<RKKYR:GfJ42/PVB9UcN,RH#D:H]]+J3P0;UP7,6S)FM4d6T\#2RNQ)AH
dL=^&Fdg5aaH]DPFCZ-#A2TcHf4/K:a@MV>=OP8-RCBX9[fF,?/U3f3UY0=\OfQJ
25]3TM27,QM63NgC;VaKG>eV:RV\b(HE(VL6CWfc,L&7SC\69Z\8+fPf<9,](9dd
ZB_6090,F]5,)b3M,&>YT:8/4]\((Bc9.V2<)D<5K[6a+fFRWO&bCTNBfKS5SVSA
,J#gB4FYOP<4X_^M/BQ<c@HF(-Q]4g^)f11#H;;E4+@^/GH-;c0?(;b#FMKMbW;V
T]W[W12&APG_<[OP1(LBGRTcc-ZXY#R@gF0PY[.6b0@:UE27a^#NGK[e(#N#5G_^
)2Fe;\IJ\JF^]5VQLNH\Uc1PC)Sb(T1cM<HH,cZSd,-\5gFLBLC-HLFZ/)c;4?(9
T_XA(EX,I^K+Q3QEYV\M[deI@AC/<V;4aM31;K_E3[[GTB7+Y6I@04V/8\c3><.G
NTSKQ,?,MGKfZKH@R@B]gX-J2H<HXS>VTE(_GJUD#fD374HL\/0(40_>X?]6\PcF
PQ8.M4cBW9>=NC/;UG8/HcDSE?(5-RP=4J7RM3-)@e3Z&g3fdUZcRE.fZUT08J0&
<bLG:?L:BC3D+5UU8Y?D.624c]LJOYc3cWA3b1OCHK=21?JS1Z8F?&<NIOC^#O>V
6LOg50ZI79\R;T8+(XG(Wb.a#Oe5&-Ma6A3GK.+Z2FAASCSYE\:.X=0T3;:>@^E;
80O?\5,G8+<^cBKJ0##/V49b@5@[D?Z/)0e@D14+4-(F-<BfL^OIF5:KQc@RJO[P
LF#[F:<gZfC1SagAVLO<dQN:9c=Y;8T)agN(V6\F.@J(/IbY)0EN@3UUdJP1fFE.
48)#d-U7A>aJ#W9NIee5G09+gcV>DI+V;/KKT:Z-PeeeS/]8)545)2EaZ.;F</J7
Z\?DWH=gC_<c3#1fL>>cF9Re(O@S9ObVZTJRg]eUPMQ/)Z&Q^-59^FGg-Y3MK,Re
);(W@RNFKDcJ=Fe1NM99&DB7SL4JgFS(^H3.\Y56U^@SDBD&E=FN<NQI4I<Rg2(?
=W<U9#>QgZDd<+O/BWQN-G^YdCO2W@?gJWdF/e_JF5)EQ4NIb_0HW48/+M1M;5gf
0d?=IPJD<]e8-Ta)dg2gRVPN=73QJIL?PB5TSc=DfI-1<H3IYK.H:;JK-7&-2R9]
D#/<>LEJ@K?=GZf1>+#X_F\H6M:<_a_8H?P,f^GW=1>R+X=^]3.1PddV@CVBV93;
aF7b2C]?=HPDLFU199+Bed7X\)XIG@L/<<9?=9H3+fc#b1H980N;e5S-VU\>IMG?
^ZIIM^P[;]fG)eOCb1O]7Q7^U_7(Bf^W)STNX5NS[UPPYACL6&V)K\HVc]D83ScA
cXJN?e6fND;MV#Y=;_F1,KKXdV\W9Z-55ZO6P:0+?WC(K5ecD?8PZ7/FBgcD3P5e
#/_730&fY3C9T#f6g8Y,W>7Na@N8c4YOS7_HcJ5Y8QUV51E](S4C4#IY__+O\1J_
.e<X@-6/\UQ#]gGFg[?B]0O.(\2Q8]NYNQgAX-Z0,?32GPC1Y\:[/&M&<bS11bZK
ecS]V)I_T/9f]-VK@_+?fMVL2F/)/JLW^J.E4MbS68L]M7S=.+QDPGe\^A?0C0<c
N6Xcc7\):F@E_d.AJ88ZdZI,.1&;][R;E<^_3d:Y@6B8O&F,9TLWF.d(_)IY86<I
PYCTd#P4c/O(EO[>=,\J)#/Y#>[1@4&SOHEeH:L9O#,b=BKZ?[\eB6PS+fD0bZO.
9^OIG?\-e[3_#Fc5gB@XWMc-f;3fe9DF?\0&LNgDHI;)A,Of[OD118]-2:K\)/c[
5KR?@agY=a&X911#=(D<>;#de-EY]I,g-d0f=\2-==CLJNaTg+:G.@;_@PCH6]RT
,g?18NaX5a8W;)31PSQ)Z(U_\>XgYCTaNZ&[Q;J21SR<#3fb(]8X/<SM:Dc@\K.(
OZ/=R2GEK0aT+:.1aHMeYNgQ,=_3ZUOCaRa8)F68b[]03[=GH,a[3dUWV)EJT>)[
)S^;8A(b;N9PQ]LH9EP-P&\W<<GX-:DY51&]gSRB2#DDZP<L2EX8>4<H3ec^G+;>
0D6I]VCR=2T\K\A#3A,2J6?04J[N.J1[^??9e+=<cb2TG&+G3-R0^UT3.L6/eL?d
PQNRRNE\B8KW1F\dM/-0T]Og-QV;JR?&IP)+C/GT4,WcTXE4+>R22W;^^E[e1XJ5
87H.S9-e);K)5OXfaIHBK6c9I0W&6:=PDTF22;7D_gMSB=E6cfN-\ZHSZ0F995=?
6DX)MWU,P6=G78NV\N7ZbAZ;d)X[.YH_>;5K8<WK6>P5b1+KY8VfLa<>_-fN>5GC
:Z1G93B##BbZYP8F\@HfP4(T4Dc2=O.D1C=3&30K6<20dXXAD(b/8^)8_gQ,ZTZ6
M>[G04C&RZ,\5THb1MYg?FZ.5eOJ/>@?]8NHfHV</0\,P;+UYfO7)5H,R[(IGRb.
?PPC2Gg/_41IO\Qg1;W<>dN3:R0Ee0]FLCZ\\D\J9?ULE(A.eRW48<#IfNT-(78d
GNb4[P1UUb?\T=?VS4<-XIHM;XC(gQU5ICE,Lc)LCG6N^RVKI931)YBTLd^S^6.4
f0Q<UJ)e6fT1EQf0B_-;(?bYGH?O[(Xe/f^L>TG=5A3JJ&[3NUA=G4,efQ=@aG+Y
cX-GX#X4#B@^.FC&P,G:a[g>Pe;&N@+d7CS4&=UcTR_EGA\,,aEF,DZ8&E20#H^3
g1P34_c.ALZSQ@e+e<BfW2,JBFffTAQFD18,#\_GbD6MK[RdTF_3/I&8Y/S\#N3^
G6-Ed].4Lb\;II56\5f/4-4&fBZbR:eKG#SG-#DR6XXgJXH<:]DI3b7ED;PHGcTM
+bH^_e-[&WO0I7H_];BB.\,Q(Sc>1LF3a9ZRA3#>T(bg?()5VZI;P^Z]e5KFJI&;
F:.(_X1S<-(3L5?#30=S8M/>5\/OYNbc0IGO(_;U^(bQa)+)H6aL\UQb7JB?a:1;
,)Agde:N^c/#^STK/gQ6FN?c8G4/Wf>7d<+H6>R(/F9]:(1F.1+)ee,D:(\8WQR9
HD3^eN6<8/&U>S.0P#)^H4R9+DJ7.cZI>]Ia/SWYYO^fYXCQ640.]WJF1E,[S)1P
BCF;[EW@H-K6&1AD<:02@BeH-;^6SGSW7FHHd]>/AKDUd^CNV;D/:J9\A6?9:Kge
fZ1Q46=^V)PBW5R),.]XR.7TIG#WgUQaN(YUG>Q8TX:g/f)U6^V.FbRZMQ6Eabfc
K?W]?F?cD55XWG2_f<3;4,I[8&HaI519#Q[]971Z<CL)_cTKb7#5O->I581OTG)9
_aF:-+e?DCg7M,^\a4+I[JR+gGXe#P.SA1P<d+2^([e_=1J58BVW=FSK?35#QJM0
:6A8(ga06Z3POAJcF^TIb=fM2g),:[a/CGe9F2YX->Z]TQ6?#>O[VYWLF+1g?.1Z
FOZ9.0F._?aK;+LGLAO/<F-^Yg[3a@e7;g,5CgT?N&gGF<OJ9GecTF&0=CGJ#aHc
#>DRUdO94C.[;[[bC=+=Y2gf9VeWYC?dZ/acCg)W8KHG4CN7<L;gfba2]/Z-^S_c
TJ9Nd2H9b)X(PV9JA2E=6)LEBC@gXRXF.P@M[A1:_-<A;]4K(R#+<;J9U\3/S&aN
#A30,KZ4E8eRQG[\eA)_01CZ_.0P:6gF@_KNF._a9EJTK2U165,&K,dMJCAR85\P
Md)S02(Z6b.4#.UJ^PbMU@QC)@,bBRb9QL:5_;&EM6?Z[WWQQ;OGR8Y1@7NbJ;XH
7fS<0Ya8HD>]aN-7SI_20RBG\QW]aP,?c9[+0:):^T&cMTO>HdQ_CKU.+7BOP#_=
+#=L6:Rb(XR@DER)D)F;f8e@PJ<0.7;,19MO/513)V2QFJ85F_F]0@KXbMc+[>X#
B7Jd-1D@RE9E7MJ3+@6c(Q8>R2SC:B[B;0&+J7QCdd,:6=&+AY>\eL752e#GD)R0
Yc6[Qab)6B@DC\]g]^+.>e:83CMJLUVBO9/4+:@=Z&c2W4#6O5D8,Xf@RaR7HM.7
166/D_7C+3P1f=@Q[.g/ZZ_W(P:O\/U8OFISH5&,Z/2HRCT>8?g>.Z:5@@PRJc#4
_6<e.WYHd8A:5S4P4U.>BZ+M0Mf@\R=IC3^TVKA1?SD)2H^C/@72^EYM10#g0(3U
/>7O,-B3ESg8-YSI>F>CX/Z[fOKWV,N&+Q)#b24>H@DZ\:YgZZW]C2Xc)^W@@S:M
>0+TeZ[O7I#fUG-Tb\3H?W?,]B.ZB@T&>6X/[F8J.NAgTO)ZTT)L#,#[+\3G\7F[
:L@bgRB4Ce#\2VSJ0PX^f7KLQGP,>.H,-&?JID(@9[HC/T&.ZNbDFH<a]K]@-6Q]
<>Ec=OU>]@36O3IU(#XN#_CbV2Jg424]TQW:SFDX)V^gV(CI=([2DHS)4)I\3(+R
.eB&-Tb;B:DA90Kf5RHUN[Q/7Mg+#SY_T.:/QfS&P0:Q5+WA/Ze(K<4\AB6O#KGI
@A=QK;(gNI-@15V<+.:SK153B<:X;d?^N?g[\//ZB_XIN;6,HHN,V01JH4P(,GT;
4F2JBZKZBINHfBP>MKgdKZ]LP0ZO]+dWT0LNBbgZBb)gGb@,+_,<AVRO:G+QLP&L
:O4&e<BCSS[.-Wa;de:#-;:,gKS=c@@YfKMecUY-W\IX2\3N+)Y7,U#WY7fb0V(C
S@VcTC+@.@Jb^<:1/CAdDIQ/4.@OI<?DCTENS=>.][0C)b]G+=aC9D^:CY(.?^d7
YW.36YL1]/@MJ&]XVb,X8V,>#C0N(6cDQ7#?>&dfO1)GX33-G^G5)Cg-P.TJX19<
T.fHQbAK>4_I[cG(9H6><W#G._NS]/:O:6UX_f\A3KYST2b\94f26VGW8V1R2;:Y
(>=4GaNZ,FdZaX//bZ0AHaMc_be@=P0_QBL(C<=bTF#b)_KS6dU#:WK3P14GB(Y5
E>,._Z&;9H[4>/g5O-:QL]N@9@X_.C>9-V6F[e0&<0DP([DS]QI]9SXQ7cfNZUXJ
6LNVYHC>=U.NQXgg\+K?]/=\9SMER[Pc20K=N4QH2c\Y^Z:U.:3BV)3;W09[c+E=
\MeR5?H>^,g@(Ob4cYC&-/#K\La#<S05Q((.:O76+TH-8^a[MT5^CX>(5f.HNNc/
>S)=Y0^YP\QT(6MWFJU.TSFdX<+=_/ZaK;IWcKDMN59M87#Uf42CX8B1N_CfT)C>
ORbDdY(D<>AM(V6CH4U3J1-W<\eYcC.1K;:fG@.BKVbRGXI.]Y3A<HgT7/faVW=/
@WTL,bAP7Fc7JT8-(>^Q\Z]ZfX-YZ\d;;/+>DPMT5^JWAU/VLdCgFS-,;QJI\dPU
G;AN,9^7+.Ef/2?@^:[IbCWXD?Rc6SI#3348(=2;6&4I,T]):WgO\YOG3S0f_U#F
E#_1XWQ9G3g=L&VRS>L&^6.\_BSECF^D7f_#IT)DL]L_?CRR=fa8ZdVY7([(,f+R
)f\/ZFObX:OC5[>AM<aYK0&+fXX7Y+PQ/3J#c[;();CZ.[ddBM6#\E4<?_Yc+(\[
4UBTg=Z3g+X#Q>6aL#GA\6^#\9H,PER-PUYG[=VDRPb/3U54eAL;_XH_6Q@7P.IQ
8I3V3TYaO.<E5Cc2K-LD#/EQJ+,E0dDHJJ7Z(Y56aWIN72#]9)Ve=;cS(7.-#X_7
-NG)+H=8cd&8[P>ZPL:Ib#1eI6fR&WE:e1,HM4e+4D5K6J\1+RHX76L#5@&N5a[Q
<L\MCV>C2GH(CVVgE&=/T/523aDLPKVEVccg1a=b/.?EO//,N_&C/++fgQGN&I0M
9I06fMGCZBZ.KUTZTN)f>MaD0c,d/HI>&X.cfD/9OQe&]FDf/W)/LU_7,;#>EF2J
(XOQf/b/7[I]CPd.?;YUBf=>Q^2Z?R:YS9cK=)-0aLO-/@7L(M6M4)IO&.&bZFZH
dDU\<(T8F3c=:49NTcUf,[<<@(@2Ub4Ye66dcWPZ)[_7(Y>[5]\6dD,MJ8QL)3N9
N60U.[BAJJ_#.OQ5gTQ/aA?a#NWZ1_]H45[KFG=D-SHEV6PM;Y41eed&,JD=G&7Y
+VN#(?\6aKMH?5Z(2FKCY?\AAM/Z7DF<()>:N+8A=A+6/70-(3XHV@?GK9c7fGSS
Z&c?VX09<)bRV>-KbgQH_\?&FP1TecO5@N/LB>7@b5JeR=UF^^EQ^QbD)F0bAQ^d
B1#P,G_c\6K-6N.G5FKJFF:T#Ee;:RYSNSP6K5_SSH<KX<<,VGcIb.JaYA?<a(cQ
W;=IZZ13VX@:66NF0(O-^<C.eSMY1K.T]5D-H/7C3VBb_:7#^_7?\=FB2cGVC:/]
bT6,XQE2L:09\2(DL?d&MR4Mb4+66)fP(AC;@FRb)UVPH.4V3(?WEK#ZSI.&+dK^
:Y<cOJ\J-f&SS6V(QMPZX)HOJ+,R-HXGP<Oe@-Gc>\E;[\@MU1E\0]6+^K0a]5PF
633UR\<(CV38_2L&Z_E:G7Z2T=/,Tf=@a=@b?WA=_POJe#C7<2ZCQ7f_T6D;Z<S<
_UGVAL-dGEeOeg6^--SX&PP>9dSJAV?>6GSS85=D(/+Y5119/^e(4C08PIZDOR7V
IYHFQAPBKM]@19&(.?PIL/RY6XU0.)O1_C)^)=AJ\^,.1@60764SSfL@NE6ZPA9&
3E1<:Q)ea]<Z^(EU@:^^DO&F5NF:,+9f<,U<@W4(1M@Mc0J<+^9HMV6.PK;QVU__
^F#];=5,80.:LVKEJ;8<aIY_]DUCC:?9UKOge,&0XCN<BZ?OW2ZSN?NR.R2;H--M
Z5df9RZ3JXg^)K=6\M?\gWS/DYWCH<HMH+>IFU]a5/0\.Y>Za(Td#+:[(R/C<75A
]/G3AUH7@\/W4WDT6;#aeM1O,7.c>9J@TYW5OYD6eg]PDFL+UJ;?^@VSa48CY;9/
H8d)^H-:)WS2<)NN04^8.+RU0d>@<+]&.AEW(T^VV7;g#2OWI+Q_dCKfV^#a&B[C
6bc3_d>a5=X50CU+L-c.FK:8.E<KFNS6@SMMN]6HE&#\9OE.5^80QUaO(?-[QG(;
@I^XW/XJPYXcS_MBN64J0>DTZFde7fIXERD202;g0JHRUb&N+1B=S4YIEfXSABf?
.:23DK^=+T/>-5c.8,I2H3@:]8F>ZN2@#AJ_e_?5G+FUV[OU>gK5+T>_GfZe>W-[
-Wc9+>ZXfPY8_51\JNFT+bNC:D2eJT>)J>PdL+,Q,\O.d#T:&F+CA[?WUeb8.C^d
[>G)cVU,/XIY/@98eWV8>LcEX=2ZX4bT9,]C5HR=//[De6AT\D>Te>;5bBf,>[D-
Q@#T=dX=IaL+;XeS\a7J+AbQf7,&0<5,f,L4YHT>c>F1)T?3+9Y-Wg<55+;V90K1
],9N75SRa5Rd8ReP2(bIC#d8AAB>&BW7g3YgV@#TR_]61PX/&9F?(P0TD:8DJV+G
cc,.UCBHbeMU0V>).)HL64<4N#.#aI:-<F1DgFMG:ECUI9)(.K(<H;0TK$
`endprotected
endmodule

module FIND_COL_TOP
`protected
0GFVL/M(^e#I(PdfEW-I5cdX[FX&ZOD->V-D[aH55N&B2fCXI5.#,)O&7->.aM9&
fWff?>EggN?A\g3D+L&cQAa+[:<3.>,O\109d)K#\54WGeRU1]I8(KUHg95[8<[5
1ORP:LIcB@K@=OPSUI.>S-9PN\V8S6Fg[#;;H+R)FT0JY<IS9gcZ(DcE>D7F5N,&
;\>ab-_+\?^DXUHR7O[/6Y091.d&Y5^3PE8B_D=Db@.TPD0;K)eV]]E)JV2>@D9c
HAGUMN5T\?(NZaA)3P9(-6.[\.PU6/7KOR(aC3.=M\feOEDV@/XQ13SP]OZ2fH@Z
(R/:Z2QP,ZQcUCJ:.;M&JRK>=bfX4cdI9HON+WP,22@X34>/Ic.-:)N>ARFW_;97
Cf,>-2Gg@RXY3E9&_+XI/V6,0QBW4aL[2/U;.fVe.W(d1#1;I->K?GbH#?<PT_;]
I&WPIDC=:gBS8L@cY2D_51:_eT(K(5WHF>C8GgL(9#^1=D7&&MdSSe?#Gc-#c=[/
,G]&_3;1LYaKK_23G5Z(XDa+/>f0+d9VW55#dB#c63d_#,[4,b9EGP50+M<.SO^/
CI45J5+K;VaCfHYHW?6WY26G&,Ig_+4bQS1#B&/MD8O^g:,=Lga-[)R=191KaWS_
N<@FC0+&><.V?#KU2J^P)?-ST<,V_WJK2fU):7RK^T#.;O/gH@gF3e2AVX[=/RRa
AI5#:_Ke7=6F>f;4=(<9/NfI(fMYN_;bE70LXab1W;S5>#:](4[_V]#f>ZEVEVP/
)F2QNc6<KNZ6,L\T/F@O9P?@-c+3P./G7^c<XR-<X9R2Ng>:A8([\Xe-&d0bWf9Q
\+>gEP2O;Z)La>?aT,]F&(+D);^&e\J9QLS7IeX9KZ^HQL+_e#]QK?1E,)N1S8P]
1]/45<-F9<5;MB<.c,DFEVSYIKPG-L1YObW-92fO3;LHE$
`endprotected
endmodule

